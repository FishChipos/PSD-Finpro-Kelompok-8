library ieee;
use ieee.std_logic_1164.all;

entity audio_equalizer is
end entity audio_equalizer;

architecture arch of audio_equalizer is
begin
end architecture arch;